//     %%%%%%%%%%%%      %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//  %%%%%%%%%%%%%%%%%%                      
// %%%%%%%%%%%%%%%%%%%% %%                
//    %% %%%%%%%%%%%%%%%%%%                
//        % %%%%%%%%%%%%%%%                 
//           %%%%%%%%%%%%%%                 ////    O P E N - S O U R C E     ////////////////////////////////////////////////////////////
//           %%%%%%%%%%%%%      %%          _________________________________////
//           %%%%%%%%%%%       %%%%                ________    _                             __      __                _     
//          %%%%%%%%%%        %%%%%%              / ____/ /_  (_)___  ____ ___  __  ______  / /__   / /   ____  ____ _(_)____ TM 
//         %%%%%%%    %%%%%%%%%%%%*%%%           / /   / __ \/ / __ \/ __ `__ \/ / / / __ \/ //_/  / /   / __ \/ __ `/ / ___/
//        %%%%% %%%%%%%%%%%%%%%%%%%%%%%         / /___/ / / / / /_/ / / / / / / /_/ / / / / ,<    / /___/ /_/ / /_/ / / /__  
//       %%%%*%%%%%%%%%%%%%  %%%%%%%%%          \____/_/ /_/_/ .___/_/ /_/ /_/\__,_/_/ /_/_/|_|  /_____/\____/\__, /_/\___/
//       %%%%%%%%%%%%%%%%%%%    %%%%%%%%%                   /_/                                              /____/  
//       %%%%%%%%%%%%%%%%                                                             ___________________________________________________               
//       %%%%%%%%%%%%%%                    //////////////////////////////////////////////       c h i p m u n k l o g i c . c o m    //// 
//         %%%%%%%%%                       
//           %%%%%%%%%%%%%%%%               
//    
//----%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//----%% 
//----%% File Name        : bram.sv
//----%% Module Name      : Dual-port Block RAM                                           
//----%% Developer        : Mitu Raj, chip@chipmunklogic.com
//----%% Vendor           : Chipmunk Logic ™ , https://chipmunklogic.com
//----%%
//----%% Description      : Simple Dual-port RAM which will be inferred on Block RAMs on FPGAs.
//----%%
//----%% Tested on        : -
//----%% Last modified on : Nov-2025
//----%% Notes            : -
//----%%                  
//----%% Copyright        : Open-source license, see README.md
//----%%                                                                                             
//----%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//###################################################################################################################################################
//                                                          D U A L - P O R T   B L O C K   R A M                                       
//###################################################################################################################################################
// Module definition
module bram #(
   // Configurable Parameters
   parameter DATA_W = 8 ,  // Data width
   parameter DEPTH  = 8 ,  // Depth

   // Derived Parameters
   parameter ADDR_W = $clog2(DEPTH) // Address width 
)(
   // Clock              
   input  logic              clk     ,   // Clock

   // Write Port
   input  logic              i_wren  ,  // Write Enable
   input  logic [ADDR_W-1:0] i_waddr ,  // Write-address                    
   input  logic [DATA_W-1:0] i_wdata ,  // Write-data 
                    
   // Read Port
   input  logic [ADDR_W-1:0] i_raddr ,  // Read-address                   
   output logic [DATA_W-1:0] o_rdata    // Read-data                   
);

// Data array
(* ram_style = "block" *)
logic [DATA_W-1:0] dt_arr_rg [DEPTH] ;

// Synchronous write
always_ff @(posedge clk) begin         
   if (i_wren) begin                          
      dt_arr_rg[i_waddr] <= i_wdata  ;      
   end
end

// Synchronous read
always_ff @(posedge clk) begin         
   o_rdata <= dt_arr_rg[i_raddr];
end

endmodule
//###################################################################################################################################################
//                                                          D U A L - P O R T   B L O C K   R A M                                       
//###################################################################################################################################################
